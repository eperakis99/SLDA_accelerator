`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input reset,
    input clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    input ap_done_reg_0,
    input ap_done_reg_1,
    input ap_done_reg_2,
    input ap_done_reg_3,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 2'b0;
    localparam ST_DL_DETECTED = 2'b1;
    localparam ST_DL_REPORT = 2'b10;

    reg find_df_deadlock = 0;
    reg [1:0] CS_fsm;
    reg [1:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg) begin
        NS_fsm = CS_fsm;
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = |dl_detect_reg;

    // dl_done_reg record the cycles has been reported
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    always @ (CS_fsm or dl_detect_reg or dl_done_reg) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_detect_reg[i] & ~dl_done_reg[i] & ~(|origin)) begin
                    origin = 'b1 << i;
                end
            end
        end
        else begin
            origin = 'b0;
        end
    end
    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [328:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "SLDA_final.Block_split2_proc_U0";
                end
                1 : begin
                    proc_path = "SLDA_final.SLDA_update_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [328:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [328:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [272:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    1: begin
                        if (~AESL_inst_SLDA_final.lambda_V_0_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_0_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_0_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_0_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_0_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_0_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_1_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_1_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_1_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_1_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_1_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_1_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_2_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_2_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_2_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_2_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_2_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_2_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_3_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_3_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_3_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_3_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_3_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_3_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_4_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_4_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_4_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_4_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_4_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_4_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_5_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_5_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_5_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_5_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_5_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_5_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_6_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_6_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_6_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_6_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_6_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_6_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_7_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_7_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_7_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_7_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_7_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_7_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_8_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_8_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_8_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_8_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_8_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_8_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_9_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_9_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_9_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_9_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_9_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_9_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_10_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_10_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_10_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_10_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_10_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_10_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_11_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_11_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_11_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_11_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_11_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_11_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_12_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_12_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_12_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_12_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_12_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_12_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_13_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_13_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_13_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_13_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_13_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_13_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_14_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_14_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_14_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_14_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_14_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_14_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_15_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_15_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_15_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_15_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_15_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_15_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_16_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_16_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_16_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_16_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_16_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_16_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_17_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_17_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_17_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_17_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_17_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_17_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_18_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_18_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_18_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_18_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_18_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_18_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_19_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_19_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_19_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_19_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_19_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_19_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_20_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_20_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_20_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_20_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_20_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_20_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_21_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_21_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_21_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_21_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_21_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_21_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_22_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_22_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_22_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_22_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_22_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_22_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_23_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_23_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_23_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_23_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_23_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_23_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_24_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_24_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_24_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_24_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_24_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_24_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_25_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_25_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_25_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_25_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_25_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_25_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_26_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_26_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_26_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_26_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_26_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_26_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_27_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_27_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_27_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_27_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_27_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_27_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_28_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_28_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_28_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_28_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_28_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_28_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_29_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_29_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_29_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_29_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_29_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_29_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_30_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_30_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_30_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_30_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_30_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_30_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_31_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_31_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_31_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_31_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_31_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_31_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_32_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_32_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_32_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_32_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_32_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_32_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_33_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_33_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_33_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_33_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_33_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_33_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_34_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_34_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_34_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_34_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_34_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_34_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_35_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_35_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_35_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_35_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_35_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_35_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_36_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_36_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_36_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_36_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_36_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_36_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_37_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_37_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_37_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_37_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_37_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_37_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_38_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_38_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_38_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_38_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_38_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_38_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_39_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_39_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_39_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_39_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_39_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_39_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_40_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_40_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_40_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_40_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_40_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_40_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_41_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_41_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_41_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_41_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_41_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_41_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_42_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_42_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_42_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_42_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_42_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_42_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_43_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_43_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_43_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_43_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_43_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_43_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_44_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_44_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_44_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_44_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_44_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_44_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_45_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_45_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_45_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_45_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_45_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_45_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_46_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_46_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_46_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_46_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_46_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_46_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_47_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_47_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_47_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_47_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_47_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_47_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_48_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_48_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_48_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_48_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_48_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_48_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_49_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_49_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_49_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_49_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_49_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_49_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_50_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_50_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_50_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_50_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_50_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_50_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_51_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_51_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_51_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_51_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_51_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_51_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_52_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_52_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_52_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_52_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_52_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_52_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_53_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_53_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_53_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_53_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_53_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_53_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_54_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_54_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_54_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_54_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_54_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_54_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_55_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_55_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_55_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_55_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_55_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_55_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_56_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_56_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_56_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_56_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_56_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_56_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_57_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_57_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_57_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_57_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_57_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_57_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_58_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_58_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_58_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_58_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_58_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_58_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_59_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_59_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_59_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_59_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_59_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_59_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_60_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_60_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_60_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_60_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_60_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_60_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_61_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_61_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_61_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_61_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_61_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_61_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_62_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_62_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_62_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_62_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_62_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_62_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_63_U.i_full_n & AESL_inst_SLDA_final.Block_split2_proc_U0.grp_init_module_fu_2804.ap_done & ap_done_reg_0 & ~AESL_inst_SLDA_final.lambda_V_63_U.t_read) begin
                            if (~AESL_inst_SLDA_final.lambda_V_63_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_63_U' written by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_63_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_63_U' read by process 'SLDA_final.SLDA_update_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (AESL_inst_SLDA_final.ap_sync_Block_split2_proc_U0_ap_ready & AESL_inst_SLDA_final.Block_split2_proc_U0.ap_idle & ~AESL_inst_SLDA_final.ap_sync_SLDA_update_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'SLDA_final.SLDA_update_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    0: begin
                        if (~AESL_inst_SLDA_final.lambda_V_0_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_0_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_0_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_0_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_0_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_0_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_1_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_1_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_1_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_1_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_1_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_1_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_10_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_10_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_10_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_10_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_10_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_10_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_10_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_10_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_11_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_11_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_11_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_11_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_11_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_11_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_11_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_11_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_12_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_12_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_12_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_12_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_12_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_12_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_12_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_12_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_13_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_13_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_13_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_13_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_13_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_13_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_13_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_13_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_14_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_14_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_14_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_14_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_14_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_14_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_14_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_14_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_15_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_15_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_15_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_15_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_15_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_15_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_15_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_15_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_16_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_16_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_16_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_16_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_16_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_16_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_16_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_16_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_17_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_17_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_17_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_17_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_17_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_17_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_17_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_17_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_18_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_18_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_18_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_18_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_18_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_18_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_18_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_18_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_19_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_19_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_19_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_19_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_19_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_19_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_19_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_19_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_2_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_2_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_2_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_2_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_2_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_2_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_20_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_20_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_20_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_20_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_20_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_20_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_20_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_20_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_21_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_21_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_21_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_21_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_21_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_21_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_21_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_21_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_22_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_22_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_22_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_22_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_22_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_22_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_22_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_22_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_23_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_23_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_23_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_23_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_23_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_23_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_23_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_23_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_24_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_24_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_24_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_24_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_24_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_24_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_24_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_24_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_25_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_25_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_25_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_25_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_25_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_25_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_25_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_25_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_26_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_26_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_26_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_26_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_26_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_26_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_26_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_26_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_27_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_27_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_27_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_27_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_27_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_27_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_27_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_27_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_28_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_28_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_28_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_28_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_28_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_28_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_28_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_28_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_29_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_29_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_29_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_29_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_29_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_29_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_29_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_29_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_3_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_3_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_3_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_3_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_3_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_3_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_30_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_30_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_30_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_30_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_30_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_30_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_30_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_30_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_31_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_31_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_31_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_31_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_31_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_31_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_31_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_31_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_32_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_32_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_32_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_32_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_32_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_32_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_32_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_32_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_33_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_33_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_33_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_33_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_33_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_33_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_33_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_33_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_34_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_34_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_34_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_34_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_34_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_34_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_34_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_34_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_35_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_35_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_35_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_35_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_35_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_35_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_35_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_35_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_36_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_36_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_36_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_36_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_36_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_36_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_36_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_36_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_37_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_37_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_37_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_37_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_37_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_37_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_37_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_37_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_38_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_38_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_38_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_38_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_38_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_38_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_38_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_38_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_39_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_39_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_39_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_39_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_39_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_39_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_39_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_39_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_4_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_4_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_4_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_4_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_4_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_4_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_40_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_40_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_40_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_40_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_40_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_40_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_40_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_40_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_41_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_41_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_41_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_41_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_41_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_41_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_41_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_41_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_42_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_42_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_42_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_42_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_42_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_42_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_42_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_42_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_43_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_43_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_43_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_43_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_43_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_43_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_43_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_43_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_44_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_44_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_44_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_44_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_44_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_44_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_44_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_44_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_45_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_45_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_45_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_45_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_45_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_45_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_45_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_45_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_46_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_46_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_46_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_46_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_46_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_46_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_46_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_46_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_47_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_47_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_47_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_47_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_47_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_47_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_47_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_47_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_48_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_48_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_48_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_48_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_48_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_48_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_48_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_48_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_49_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_49_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_49_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_49_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_49_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_49_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_49_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_49_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_5_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_5_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_5_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_5_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_5_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_5_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_50_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_50_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_50_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_50_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_50_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_50_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_50_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_50_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_51_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_51_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_51_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_51_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_51_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_51_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_51_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_51_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_52_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_52_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_52_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_52_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_52_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_52_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_52_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_52_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_53_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_53_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_53_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_53_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_53_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_53_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_53_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_53_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_54_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_54_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_54_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_54_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_54_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_54_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_54_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_54_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_55_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_55_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_55_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_55_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_55_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_55_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_55_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_55_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_56_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_56_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_56_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_56_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_56_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_56_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_56_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_56_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_57_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_57_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_57_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_57_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_57_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_57_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_57_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_57_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_58_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_58_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_58_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_58_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_58_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_58_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_58_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_58_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_59_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_59_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_59_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_59_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_59_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_59_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_59_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_59_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_6_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_6_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_6_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_6_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_6_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_6_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_60_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_60_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_60_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_60_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_60_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_60_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_60_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_60_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_61_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_61_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_61_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_61_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_61_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_61_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_61_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_61_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_62_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_62_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_62_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_62_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_62_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_62_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_62_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_62_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_63_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_63_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_63_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_63_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_63_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_63_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_63_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_63_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_7_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_7_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_7_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_7_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_7_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_7_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_7_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_7_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_8_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_8_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_8_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_8_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_8_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_8_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_8_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_8_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~AESL_inst_SLDA_final.lambda_V_9_U.t_empty_n & AESL_inst_SLDA_final.SLDA_update_U0.grp_compute_weights_with_matrix_mult_fu_1604.ap_idle & ~AESL_inst_SLDA_final.lambda_V_9_U.i_write) begin
                            if (~AESL_inst_SLDA_final.lambda_V_9_U.t_empty_n) begin
                                $display("//      Blocked by empty input PIPO 'SLDA_final.lambda_V_9_U' written by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_9_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_SLDA_final.lambda_V_9_U.i_full_n) begin
                                $display("//      Blocked by full output PIPO 'SLDA_final.lambda_V_9_U' read by process 'SLDA_final.Block_split2_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path SLDA_final.lambda_V_9_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (AESL_inst_SLDA_final.ap_sync_SLDA_update_U0_ap_ready & AESL_inst_SLDA_final.SLDA_update_U0.ap_idle & ~AESL_inst_SLDA_final.ap_sync_Block_split2_proc_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'SLDA_final.Block_split2_proc_U0'");
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        find_df_deadlock = 1;
                        @(negedge clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
